mypll_inst: mypll
port map(
          PACKAGEPIN => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => ,
          BYPASS => ,
          LOCK => 
        );
