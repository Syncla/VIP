// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jan 19 2018 14:26:32

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Blink" view "INTERFACE"

module Blink (
    ref_clk,
    led,
    clk);

    input ref_clk;
    output led;
    output clk;

    wire N__1486;
    wire N__1472;
    wire N__1471;
    wire N__1470;
    wire N__1463;
    wire N__1462;
    wire N__1461;
    wire N__1444;
    wire N__1443;
    wire N__1442;
    wire N__1441;
    wire N__1438;
    wire N__1433;
    wire N__1430;
    wire N__1427;
    wire N__1420;
    wire N__1419;
    wire N__1418;
    wire N__1417;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1399;
    wire N__1396;
    wire N__1393;
    wire N__1390;
    wire N__1389;
    wire N__1388;
    wire N__1387;
    wire N__1386;
    wire N__1385;
    wire N__1378;
    wire N__1371;
    wire N__1366;
    wire N__1365;
    wire N__1364;
    wire N__1363;
    wire N__1362;
    wire N__1359;
    wire N__1356;
    wire N__1353;
    wire N__1344;
    wire N__1339;
    wire N__1336;
    wire N__1333;
    wire N__1332;
    wire N__1329;
    wire N__1326;
    wire N__1321;
    wire N__1320;
    wire N__1317;
    wire N__1314;
    wire N__1309;
    wire N__1308;
    wire N__1305;
    wire N__1302;
    wire N__1297;
    wire N__1296;
    wire N__1291;
    wire N__1288;
    wire N__1287;
    wire N__1286;
    wire N__1285;
    wire N__1278;
    wire N__1277;
    wire N__1274;
    wire N__1271;
    wire N__1268;
    wire N__1261;
    wire N__1260;
    wire N__1259;
    wire N__1258;
    wire N__1257;
    wire N__1256;
    wire N__1255;
    wire N__1254;
    wire N__1253;
    wire N__1252;
    wire N__1243;
    wire N__1240;
    wire N__1231;
    wire N__1228;
    wire N__1225;
    wire N__1216;
    wire N__1215;
    wire N__1214;
    wire N__1213;
    wire N__1210;
    wire N__1207;
    wire N__1204;
    wire N__1201;
    wire N__1196;
    wire N__1193;
    wire N__1186;
    wire N__1183;
    wire N__1182;
    wire N__1179;
    wire N__1176;
    wire N__1173;
    wire N__1170;
    wire N__1165;
    wire N__1162;
    wire N__1161;
    wire N__1158;
    wire N__1157;
    wire N__1156;
    wire N__1155;
    wire N__1154;
    wire N__1153;
    wire N__1152;
    wire N__1135;
    wire N__1132;
    wire N__1129;
    wire N__1126;
    wire N__1125;
    wire N__1124;
    wire N__1123;
    wire N__1120;
    wire N__1117;
    wire N__1114;
    wire N__1111;
    wire N__1102;
    wire N__1101;
    wire N__1100;
    wire N__1099;
    wire N__1096;
    wire N__1093;
    wire N__1090;
    wire N__1087;
    wire N__1078;
    wire N__1077;
    wire N__1076;
    wire N__1073;
    wire N__1070;
    wire N__1067;
    wire N__1066;
    wire N__1063;
    wire N__1058;
    wire N__1055;
    wire N__1048;
    wire N__1047;
    wire N__1046;
    wire N__1045;
    wire N__1042;
    wire N__1039;
    wire N__1036;
    wire N__1033;
    wire N__1024;
    wire N__1021;
    wire N__1018;
    wire N__1015;
    wire N__1012;
    wire N__1009;
    wire N__1006;
    wire N__1003;
    wire N__1000;
    wire N__997;
    wire N__994;
    wire N__991;
    wire N__988;
    wire N__985;
    wire N__982;
    wire N__981;
    wire N__976;
    wire N__973;
    wire N__970;
    wire N__967;
    wire N__964;
    wire N__963;
    wire N__962;
    wire N__961;
    wire N__954;
    wire N__951;
    wire N__946;
    wire N__943;
    wire N__942;
    wire N__941;
    wire N__940;
    wire N__933;
    wire N__930;
    wire N__925;
    wire N__922;
    wire N__919;
    wire N__916;
    wire N__913;
    wire N__910;
    wire N__907;
    wire N__904;
    wire N__903;
    wire N__900;
    wire N__897;
    wire N__892;
    wire N__889;
    wire N__886;
    wire N__885;
    wire N__882;
    wire N__879;
    wire N__874;
    wire N__873;
    wire N__870;
    wire N__867;
    wire N__862;
    wire N__859;
    wire N__858;
    wire N__855;
    wire N__852;
    wire N__847;
    wire N__846;
    wire N__843;
    wire N__840;
    wire N__835;
    wire N__834;
    wire N__831;
    wire N__828;
    wire N__823;
    wire N__820;
    wire N__819;
    wire N__816;
    wire N__813;
    wire N__808;
    wire N__805;
    wire N__802;
    wire N__801;
    wire N__800;
    wire N__797;
    wire N__792;
    wire N__789;
    wire N__784;
    wire N__781;
    wire N__778;
    wire N__777;
    wire N__774;
    wire N__771;
    wire N__768;
    wire N__763;
    wire N__760;
    wire N__757;
    wire N__754;
    wire N__751;
    wire N__748;
    wire N__745;
    wire N__742;
    wire N__739;
    wire N__736;
    wire N__733;
    wire N__730;
    wire N__727;
    wire N__724;
    wire N__721;
    wire N__718;
    wire N__715;
    wire N__712;
    wire N__709;
    wire N__706;
    wire N__703;
    wire N__700;
    wire N__697;
    wire N__694;
    wire N__691;
    wire N__688;
    wire N__685;
    wire N__682;
    wire N__679;
    wire N__676;
    wire N__673;
    wire N__670;
    wire N__667;
    wire N__664;
    wire \mypll_inst.clk_c ;
    wire VCCG0;
    wire GNDG0;
    wire GB_BUFFER_clk_c_g_THRU_CO;
    wire bfn_7_1_0_;
    wire countZ0Z_2;
    wire un2_count_1_cry_1;
    wire countZ0Z_3;
    wire un2_count_1_cry_2;
    wire countZ0Z_4;
    wire un2_count_1_cry_3;
    wire un2_count_1_cry_4;
    wire un2_count_1_cry_5;
    wire un2_count_1_cry_6;
    wire un2_count_1_cry_7;
    wire un2_count_1_cry_8;
    wire bfn_7_2_0_;
    wire un2_count_1_cry_9;
    wire un2_count_1_cry_10;
    wire un2_count_1_cry_11;
    wire un2_count_1_cry_12;
    wire un2_count_1_cry_13;
    wire un2_count_1_cry_14;
    wire un2_count_1_cry_15;
    wire un2_count_1_cry_16;
    wire bfn_7_3_0_;
    wire un2_count_1_cry_17;
    wire un2_count_1_cry_18;
    wire un2_count_1_cry_19;
    wire un2_count_1_cry_20;
    wire un2_count_1_cry_21;
    wire count_RNO_0Z0Z_7;
    wire countZ0Z_1;
    wire count_RNO_0Z0Z_5;
    wire countZ0Z_9;
    wire countZ0Z_8;
    wire countZ0Z_10;
    wire countZ0Z_11;
    wire countZ0Z_7;
    wire op_lt_op_lt_count8lto11_2_cascade_;
    wire countZ0Z_5;
    wire op_lt_op_lt_count8lt14_cascade_;
    wire op_lt_op_lt_count8lto19_1_N_5_cascade_;
    wire countZ0Z_0;
    wire count_RNO_0Z0Z_6;
    wire countZ0Z_6;
    wire op_lt_op_lt_count8lto22_2_0_tz_cascade_;
    wire count_RNO_0Z0Z_22;
    wire count_RNO_0Z0Z_13;
    wire op_lt_op_lt_count8lto22_cascade_;
    wire op_lt_op_lt_count8lto14_0_0_cascade_;
    wire op_lt_op_lt_count8lt14;
    wire count_RNO_0Z0Z_12;
    wire op_lt_op_lt_count8lt17_cascade_;
    wire countZ0Z_16;
    wire countZ0Z_15;
    wire count_RNO_0Z0Z_21;
    wire count_RNO_0Z0Z_17;
    wire countZ0Z_18;
    wire countZ0Z_19;
    wire count_RNO_0Z0Z_14;
    wire op_lt_op_lt_count8lto19_0_cascade_;
    wire op_lt_op_lt_count8lto19_0;
    wire op_lt_op_lt_count8lt17;
    wire count_RNO_0Z0Z_20;
    wire countZ0Z_22;
    wire countZ0Z_21;
    wire countZ0Z_20;
    wire op_lt_op_lt_count8lto22_1;
    wire op_lt_op_lt_count8lto19_1_m4_i_a3_0;
    wire op_lt_op_lt_count8lto22;
    wire op_lt_op_lt_count8lto19_1_N_5;
    wire led_c;
    wire clk_c_g;
    wire countZ0Z_14;
    wire countZ0Z_13;
    wire countZ0Z_17;
    wire countZ0Z_12;
    wire op_lt_op_lt_count8lto22_d_a0_1;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \mypll_inst.mypll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \mypll_inst.mypll_inst_pll .TEST_MODE=1'b0;
    defparam \mypll_inst.mypll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \mypll_inst.mypll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \mypll_inst.mypll_inst_pll .FILTER_RANGE=3'b001;
    defparam \mypll_inst.mypll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \mypll_inst.mypll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \mypll_inst.mypll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \mypll_inst.mypll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \mypll_inst.mypll_inst_pll .DIVR=4'b0000;
    defparam \mypll_inst.mypll_inst_pll .DIVQ=3'b100;
    defparam \mypll_inst.mypll_inst_pll .DIVF=7'b0111111;
    defparam \mypll_inst.mypll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \mypll_inst.mypll_inst_pll  (
            .PLLOUTGLOBAL(),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__1018),
            .PLLOUTCORE(\mypll_inst.clk_c ),
            .LOCK(),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__1486));
    IO_PAD \mypll_inst.mypll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__1486),
            .PACKAGEPIN(ref_clk));
    IO_PAD led_obuf_iopad (
            .OE(N__1472),
            .DIN(N__1471),
            .DOUT(N__1470),
            .PACKAGEPIN(led));
    defparam led_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_preio (
            .PADOEN(N__1472),
            .PADOUT(N__1471),
            .PADIN(N__1470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_obuf_iopad (
            .OE(N__1463),
            .DIN(N__1462),
            .DOUT(N__1461),
            .PACKAGEPIN(clk));
    defparam clk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clk_obuf_preio (
            .PADOEN(N__1463),
            .PADOUT(N__1462),
            .PADIN(N__1461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__694),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__318 (
            .O(N__1444),
            .I(N__1438));
    InMux I__317 (
            .O(N__1443),
            .I(N__1433));
    InMux I__316 (
            .O(N__1442),
            .I(N__1433));
    InMux I__315 (
            .O(N__1441),
            .I(N__1430));
    InMux I__314 (
            .O(N__1438),
            .I(N__1427));
    LocalMux I__313 (
            .O(N__1433),
            .I(countZ0Z_18));
    LocalMux I__312 (
            .O(N__1430),
            .I(countZ0Z_18));
    LocalMux I__311 (
            .O(N__1427),
            .I(countZ0Z_18));
    InMux I__310 (
            .O(N__1420),
            .I(N__1412));
    InMux I__309 (
            .O(N__1419),
            .I(N__1412));
    InMux I__308 (
            .O(N__1418),
            .I(N__1409));
    InMux I__307 (
            .O(N__1417),
            .I(N__1406));
    LocalMux I__306 (
            .O(N__1412),
            .I(countZ0Z_19));
    LocalMux I__305 (
            .O(N__1409),
            .I(countZ0Z_19));
    LocalMux I__304 (
            .O(N__1406),
            .I(countZ0Z_19));
    InMux I__303 (
            .O(N__1399),
            .I(N__1396));
    LocalMux I__302 (
            .O(N__1396),
            .I(count_RNO_0Z0Z_14));
    CascadeMux I__301 (
            .O(N__1393),
            .I(op_lt_op_lt_count8lto19_0_cascade_));
    InMux I__300 (
            .O(N__1390),
            .I(N__1378));
    InMux I__299 (
            .O(N__1389),
            .I(N__1378));
    InMux I__298 (
            .O(N__1388),
            .I(N__1378));
    InMux I__297 (
            .O(N__1387),
            .I(N__1371));
    InMux I__296 (
            .O(N__1386),
            .I(N__1371));
    InMux I__295 (
            .O(N__1385),
            .I(N__1371));
    LocalMux I__294 (
            .O(N__1378),
            .I(op_lt_op_lt_count8lto19_0));
    LocalMux I__293 (
            .O(N__1371),
            .I(op_lt_op_lt_count8lto19_0));
    CascadeMux I__292 (
            .O(N__1366),
            .I(N__1359));
    CascadeMux I__291 (
            .O(N__1365),
            .I(N__1356));
    InMux I__290 (
            .O(N__1364),
            .I(N__1353));
    InMux I__289 (
            .O(N__1363),
            .I(N__1344));
    InMux I__288 (
            .O(N__1362),
            .I(N__1344));
    InMux I__287 (
            .O(N__1359),
            .I(N__1344));
    InMux I__286 (
            .O(N__1356),
            .I(N__1344));
    LocalMux I__285 (
            .O(N__1353),
            .I(op_lt_op_lt_count8lt17));
    LocalMux I__284 (
            .O(N__1344),
            .I(op_lt_op_lt_count8lt17));
    InMux I__283 (
            .O(N__1339),
            .I(N__1336));
    LocalMux I__282 (
            .O(N__1336),
            .I(count_RNO_0Z0Z_20));
    InMux I__281 (
            .O(N__1333),
            .I(N__1329));
    InMux I__280 (
            .O(N__1332),
            .I(N__1326));
    LocalMux I__279 (
            .O(N__1329),
            .I(countZ0Z_22));
    LocalMux I__278 (
            .O(N__1326),
            .I(countZ0Z_22));
    InMux I__277 (
            .O(N__1321),
            .I(N__1317));
    InMux I__276 (
            .O(N__1320),
            .I(N__1314));
    LocalMux I__275 (
            .O(N__1317),
            .I(countZ0Z_21));
    LocalMux I__274 (
            .O(N__1314),
            .I(countZ0Z_21));
    InMux I__273 (
            .O(N__1309),
            .I(N__1305));
    InMux I__272 (
            .O(N__1308),
            .I(N__1302));
    LocalMux I__271 (
            .O(N__1305),
            .I(countZ0Z_20));
    LocalMux I__270 (
            .O(N__1302),
            .I(countZ0Z_20));
    InMux I__269 (
            .O(N__1297),
            .I(N__1291));
    InMux I__268 (
            .O(N__1296),
            .I(N__1291));
    LocalMux I__267 (
            .O(N__1291),
            .I(op_lt_op_lt_count8lto22_1));
    InMux I__266 (
            .O(N__1288),
            .I(N__1278));
    InMux I__265 (
            .O(N__1287),
            .I(N__1278));
    InMux I__264 (
            .O(N__1286),
            .I(N__1278));
    InMux I__263 (
            .O(N__1285),
            .I(N__1274));
    LocalMux I__262 (
            .O(N__1278),
            .I(N__1271));
    InMux I__261 (
            .O(N__1277),
            .I(N__1268));
    LocalMux I__260 (
            .O(N__1274),
            .I(op_lt_op_lt_count8lto19_1_m4_i_a3_0));
    Odrv4 I__259 (
            .O(N__1271),
            .I(op_lt_op_lt_count8lto19_1_m4_i_a3_0));
    LocalMux I__258 (
            .O(N__1268),
            .I(op_lt_op_lt_count8lto19_1_m4_i_a3_0));
    InMux I__257 (
            .O(N__1261),
            .I(N__1243));
    InMux I__256 (
            .O(N__1260),
            .I(N__1243));
    InMux I__255 (
            .O(N__1259),
            .I(N__1243));
    InMux I__254 (
            .O(N__1258),
            .I(N__1243));
    InMux I__253 (
            .O(N__1257),
            .I(N__1240));
    InMux I__252 (
            .O(N__1256),
            .I(N__1231));
    InMux I__251 (
            .O(N__1255),
            .I(N__1231));
    InMux I__250 (
            .O(N__1254),
            .I(N__1231));
    InMux I__249 (
            .O(N__1253),
            .I(N__1231));
    InMux I__248 (
            .O(N__1252),
            .I(N__1228));
    LocalMux I__247 (
            .O(N__1243),
            .I(N__1225));
    LocalMux I__246 (
            .O(N__1240),
            .I(op_lt_op_lt_count8lto22));
    LocalMux I__245 (
            .O(N__1231),
            .I(op_lt_op_lt_count8lto22));
    LocalMux I__244 (
            .O(N__1228),
            .I(op_lt_op_lt_count8lto22));
    Odrv4 I__243 (
            .O(N__1225),
            .I(op_lt_op_lt_count8lto22));
    CascadeMux I__242 (
            .O(N__1216),
            .I(N__1210));
    CascadeMux I__241 (
            .O(N__1215),
            .I(N__1207));
    CascadeMux I__240 (
            .O(N__1214),
            .I(N__1204));
    InMux I__239 (
            .O(N__1213),
            .I(N__1201));
    InMux I__238 (
            .O(N__1210),
            .I(N__1196));
    InMux I__237 (
            .O(N__1207),
            .I(N__1196));
    InMux I__236 (
            .O(N__1204),
            .I(N__1193));
    LocalMux I__235 (
            .O(N__1201),
            .I(op_lt_op_lt_count8lto19_1_N_5));
    LocalMux I__234 (
            .O(N__1196),
            .I(op_lt_op_lt_count8lto19_1_N_5));
    LocalMux I__233 (
            .O(N__1193),
            .I(op_lt_op_lt_count8lto19_1_N_5));
    IoInMux I__232 (
            .O(N__1186),
            .I(N__1183));
    LocalMux I__231 (
            .O(N__1183),
            .I(N__1179));
    CascadeMux I__230 (
            .O(N__1182),
            .I(N__1176));
    Span4Mux_s0_v I__229 (
            .O(N__1179),
            .I(N__1173));
    InMux I__228 (
            .O(N__1176),
            .I(N__1170));
    Odrv4 I__227 (
            .O(N__1173),
            .I(led_c));
    LocalMux I__226 (
            .O(N__1170),
            .I(led_c));
    InMux I__225 (
            .O(N__1165),
            .I(N__1162));
    LocalMux I__224 (
            .O(N__1162),
            .I(N__1158));
    ClkMux I__223 (
            .O(N__1161),
            .I(N__1135));
    Glb2LocalMux I__222 (
            .O(N__1158),
            .I(N__1135));
    ClkMux I__221 (
            .O(N__1157),
            .I(N__1135));
    ClkMux I__220 (
            .O(N__1156),
            .I(N__1135));
    ClkMux I__219 (
            .O(N__1155),
            .I(N__1135));
    ClkMux I__218 (
            .O(N__1154),
            .I(N__1135));
    ClkMux I__217 (
            .O(N__1153),
            .I(N__1135));
    ClkMux I__216 (
            .O(N__1152),
            .I(N__1135));
    GlobalMux I__215 (
            .O(N__1135),
            .I(N__1132));
    gio2CtrlBuf I__214 (
            .O(N__1132),
            .I(clk_c_g));
    InMux I__213 (
            .O(N__1129),
            .I(N__1126));
    LocalMux I__212 (
            .O(N__1126),
            .I(N__1120));
    InMux I__211 (
            .O(N__1125),
            .I(N__1117));
    InMux I__210 (
            .O(N__1124),
            .I(N__1114));
    InMux I__209 (
            .O(N__1123),
            .I(N__1111));
    Odrv4 I__208 (
            .O(N__1120),
            .I(countZ0Z_14));
    LocalMux I__207 (
            .O(N__1117),
            .I(countZ0Z_14));
    LocalMux I__206 (
            .O(N__1114),
            .I(countZ0Z_14));
    LocalMux I__205 (
            .O(N__1111),
            .I(countZ0Z_14));
    InMux I__204 (
            .O(N__1102),
            .I(N__1096));
    InMux I__203 (
            .O(N__1101),
            .I(N__1093));
    InMux I__202 (
            .O(N__1100),
            .I(N__1090));
    InMux I__201 (
            .O(N__1099),
            .I(N__1087));
    LocalMux I__200 (
            .O(N__1096),
            .I(countZ0Z_13));
    LocalMux I__199 (
            .O(N__1093),
            .I(countZ0Z_13));
    LocalMux I__198 (
            .O(N__1090),
            .I(countZ0Z_13));
    LocalMux I__197 (
            .O(N__1087),
            .I(countZ0Z_13));
    CascadeMux I__196 (
            .O(N__1078),
            .I(N__1073));
    CascadeMux I__195 (
            .O(N__1077),
            .I(N__1070));
    CascadeMux I__194 (
            .O(N__1076),
            .I(N__1067));
    InMux I__193 (
            .O(N__1073),
            .I(N__1063));
    InMux I__192 (
            .O(N__1070),
            .I(N__1058));
    InMux I__191 (
            .O(N__1067),
            .I(N__1058));
    InMux I__190 (
            .O(N__1066),
            .I(N__1055));
    LocalMux I__189 (
            .O(N__1063),
            .I(countZ0Z_17));
    LocalMux I__188 (
            .O(N__1058),
            .I(countZ0Z_17));
    LocalMux I__187 (
            .O(N__1055),
            .I(countZ0Z_17));
    InMux I__186 (
            .O(N__1048),
            .I(N__1042));
    InMux I__185 (
            .O(N__1047),
            .I(N__1039));
    InMux I__184 (
            .O(N__1046),
            .I(N__1036));
    InMux I__183 (
            .O(N__1045),
            .I(N__1033));
    LocalMux I__182 (
            .O(N__1042),
            .I(countZ0Z_12));
    LocalMux I__181 (
            .O(N__1039),
            .I(countZ0Z_12));
    LocalMux I__180 (
            .O(N__1036),
            .I(countZ0Z_12));
    LocalMux I__179 (
            .O(N__1033),
            .I(countZ0Z_12));
    InMux I__178 (
            .O(N__1024),
            .I(N__1021));
    LocalMux I__177 (
            .O(N__1021),
            .I(op_lt_op_lt_count8lto22_d_a0_1));
    IoInMux I__176 (
            .O(N__1018),
            .I(N__1015));
    LocalMux I__175 (
            .O(N__1015),
            .I(N__1012));
    Span4Mux_s0_v I__174 (
            .O(N__1012),
            .I(N__1009));
    Odrv4 I__173 (
            .O(N__1009),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__172 (
            .O(N__1006),
            .I(op_lt_op_lt_count8lto22_2_0_tz_cascade_));
    InMux I__171 (
            .O(N__1003),
            .I(N__1000));
    LocalMux I__170 (
            .O(N__1000),
            .I(count_RNO_0Z0Z_22));
    InMux I__169 (
            .O(N__997),
            .I(N__994));
    LocalMux I__168 (
            .O(N__994),
            .I(N__991));
    Odrv4 I__167 (
            .O(N__991),
            .I(count_RNO_0Z0Z_13));
    CascadeMux I__166 (
            .O(N__988),
            .I(op_lt_op_lt_count8lto22_cascade_));
    CascadeMux I__165 (
            .O(N__985),
            .I(op_lt_op_lt_count8lto14_0_0_cascade_));
    InMux I__164 (
            .O(N__982),
            .I(N__976));
    InMux I__163 (
            .O(N__981),
            .I(N__976));
    LocalMux I__162 (
            .O(N__976),
            .I(op_lt_op_lt_count8lt14));
    InMux I__161 (
            .O(N__973),
            .I(N__970));
    LocalMux I__160 (
            .O(N__970),
            .I(count_RNO_0Z0Z_12));
    CascadeMux I__159 (
            .O(N__967),
            .I(op_lt_op_lt_count8lt17_cascade_));
    InMux I__158 (
            .O(N__964),
            .I(N__954));
    InMux I__157 (
            .O(N__963),
            .I(N__954));
    InMux I__156 (
            .O(N__962),
            .I(N__954));
    InMux I__155 (
            .O(N__961),
            .I(N__951));
    LocalMux I__154 (
            .O(N__954),
            .I(countZ0Z_16));
    LocalMux I__153 (
            .O(N__951),
            .I(countZ0Z_16));
    CascadeMux I__152 (
            .O(N__946),
            .I(N__943));
    InMux I__151 (
            .O(N__943),
            .I(N__933));
    InMux I__150 (
            .O(N__942),
            .I(N__933));
    InMux I__149 (
            .O(N__941),
            .I(N__933));
    InMux I__148 (
            .O(N__940),
            .I(N__930));
    LocalMux I__147 (
            .O(N__933),
            .I(countZ0Z_15));
    LocalMux I__146 (
            .O(N__930),
            .I(countZ0Z_15));
    InMux I__145 (
            .O(N__925),
            .I(N__922));
    LocalMux I__144 (
            .O(N__922),
            .I(count_RNO_0Z0Z_21));
    CascadeMux I__143 (
            .O(N__919),
            .I(N__916));
    InMux I__142 (
            .O(N__916),
            .I(N__913));
    LocalMux I__141 (
            .O(N__913),
            .I(count_RNO_0Z0Z_17));
    InMux I__140 (
            .O(N__910),
            .I(N__907));
    LocalMux I__139 (
            .O(N__907),
            .I(count_RNO_0Z0Z_7));
    InMux I__138 (
            .O(N__904),
            .I(N__900));
    InMux I__137 (
            .O(N__903),
            .I(N__897));
    LocalMux I__136 (
            .O(N__900),
            .I(countZ0Z_1));
    LocalMux I__135 (
            .O(N__897),
            .I(countZ0Z_1));
    InMux I__134 (
            .O(N__892),
            .I(N__889));
    LocalMux I__133 (
            .O(N__889),
            .I(count_RNO_0Z0Z_5));
    InMux I__132 (
            .O(N__886),
            .I(N__882));
    InMux I__131 (
            .O(N__885),
            .I(N__879));
    LocalMux I__130 (
            .O(N__882),
            .I(countZ0Z_9));
    LocalMux I__129 (
            .O(N__879),
            .I(countZ0Z_9));
    InMux I__128 (
            .O(N__874),
            .I(N__870));
    InMux I__127 (
            .O(N__873),
            .I(N__867));
    LocalMux I__126 (
            .O(N__870),
            .I(countZ0Z_8));
    LocalMux I__125 (
            .O(N__867),
            .I(countZ0Z_8));
    CascadeMux I__124 (
            .O(N__862),
            .I(N__859));
    InMux I__123 (
            .O(N__859),
            .I(N__855));
    InMux I__122 (
            .O(N__858),
            .I(N__852));
    LocalMux I__121 (
            .O(N__855),
            .I(countZ0Z_10));
    LocalMux I__120 (
            .O(N__852),
            .I(countZ0Z_10));
    InMux I__119 (
            .O(N__847),
            .I(N__843));
    InMux I__118 (
            .O(N__846),
            .I(N__840));
    LocalMux I__117 (
            .O(N__843),
            .I(countZ0Z_11));
    LocalMux I__116 (
            .O(N__840),
            .I(countZ0Z_11));
    InMux I__115 (
            .O(N__835),
            .I(N__831));
    InMux I__114 (
            .O(N__834),
            .I(N__828));
    LocalMux I__113 (
            .O(N__831),
            .I(countZ0Z_7));
    LocalMux I__112 (
            .O(N__828),
            .I(countZ0Z_7));
    CascadeMux I__111 (
            .O(N__823),
            .I(op_lt_op_lt_count8lto11_2_cascade_));
    InMux I__110 (
            .O(N__820),
            .I(N__816));
    InMux I__109 (
            .O(N__819),
            .I(N__813));
    LocalMux I__108 (
            .O(N__816),
            .I(countZ0Z_5));
    LocalMux I__107 (
            .O(N__813),
            .I(countZ0Z_5));
    CascadeMux I__106 (
            .O(N__808),
            .I(op_lt_op_lt_count8lt14_cascade_));
    CascadeMux I__105 (
            .O(N__805),
            .I(op_lt_op_lt_count8lto19_1_N_5_cascade_));
    CascadeMux I__104 (
            .O(N__802),
            .I(N__797));
    InMux I__103 (
            .O(N__801),
            .I(N__792));
    InMux I__102 (
            .O(N__800),
            .I(N__792));
    InMux I__101 (
            .O(N__797),
            .I(N__789));
    LocalMux I__100 (
            .O(N__792),
            .I(countZ0Z_0));
    LocalMux I__99 (
            .O(N__789),
            .I(countZ0Z_0));
    InMux I__98 (
            .O(N__784),
            .I(N__781));
    LocalMux I__97 (
            .O(N__781),
            .I(count_RNO_0Z0Z_6));
    CascadeMux I__96 (
            .O(N__778),
            .I(N__774));
    InMux I__95 (
            .O(N__777),
            .I(N__771));
    InMux I__94 (
            .O(N__774),
            .I(N__768));
    LocalMux I__93 (
            .O(N__771),
            .I(countZ0Z_6));
    LocalMux I__92 (
            .O(N__768),
            .I(countZ0Z_6));
    InMux I__91 (
            .O(N__763),
            .I(un2_count_1_cry_13));
    InMux I__90 (
            .O(N__760),
            .I(un2_count_1_cry_14));
    InMux I__89 (
            .O(N__757),
            .I(un2_count_1_cry_15));
    InMux I__88 (
            .O(N__754),
            .I(bfn_7_3_0_));
    InMux I__87 (
            .O(N__751),
            .I(un2_count_1_cry_17));
    InMux I__86 (
            .O(N__748),
            .I(un2_count_1_cry_18));
    InMux I__85 (
            .O(N__745),
            .I(un2_count_1_cry_19));
    InMux I__84 (
            .O(N__742),
            .I(un2_count_1_cry_20));
    InMux I__83 (
            .O(N__739),
            .I(un2_count_1_cry_21));
    InMux I__82 (
            .O(N__736),
            .I(un2_count_1_cry_4));
    InMux I__81 (
            .O(N__733),
            .I(un2_count_1_cry_5));
    InMux I__80 (
            .O(N__730),
            .I(un2_count_1_cry_6));
    InMux I__79 (
            .O(N__727),
            .I(un2_count_1_cry_7));
    InMux I__78 (
            .O(N__724),
            .I(bfn_7_2_0_));
    InMux I__77 (
            .O(N__721),
            .I(un2_count_1_cry_9));
    InMux I__76 (
            .O(N__718),
            .I(un2_count_1_cry_10));
    InMux I__75 (
            .O(N__715),
            .I(un2_count_1_cry_11));
    InMux I__74 (
            .O(N__712),
            .I(un2_count_1_cry_12));
    IoInMux I__73 (
            .O(N__709),
            .I(N__706));
    LocalMux I__72 (
            .O(N__706),
            .I(N__703));
    Span12Mux_s8_v I__71 (
            .O(N__703),
            .I(N__700));
    Span12Mux_v I__70 (
            .O(N__700),
            .I(N__697));
    Odrv12 I__69 (
            .O(N__697),
            .I(\mypll_inst.clk_c ));
    IoInMux I__68 (
            .O(N__694),
            .I(N__691));
    LocalMux I__67 (
            .O(N__691),
            .I(GB_BUFFER_clk_c_g_THRU_CO));
    InMux I__66 (
            .O(N__688),
            .I(N__685));
    LocalMux I__65 (
            .O(N__685),
            .I(countZ0Z_2));
    InMux I__64 (
            .O(N__682),
            .I(un2_count_1_cry_1));
    InMux I__63 (
            .O(N__679),
            .I(N__676));
    LocalMux I__62 (
            .O(N__676),
            .I(countZ0Z_3));
    InMux I__61 (
            .O(N__673),
            .I(un2_count_1_cry_2));
    InMux I__60 (
            .O(N__670),
            .I(N__667));
    LocalMux I__59 (
            .O(N__667),
            .I(countZ0Z_4));
    InMux I__58 (
            .O(N__664),
            .I(un2_count_1_cry_3));
    defparam IN_MUX_bfv_7_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_1_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(un2_count_1_cry_8),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(un2_count_1_cry_16),
            .carryinitout(bfn_7_3_0_));
    ICE_GB \mypll_inst.PLLOUTCORE_derived_clock_RNIF7IB  (
            .USERSIGNALTOGLOBALBUFFER(N__709),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam GB_BUFFER_clk_c_g_THRU_LUT4_0_LC_5_1_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_c_g_THRU_LUT4_0_LC_5_1_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_c_g_THRU_LUT4_0_LC_5_1_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_c_g_THRU_LUT4_0_LC_5_1_6 (
            .in0(N__1165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_count_1_cry_1_c_LC_7_1_0.C_ON=1'b1;
    defparam un2_count_1_cry_1_c_LC_7_1_0.SEQ_MODE=4'b0000;
    defparam un2_count_1_cry_1_c_LC_7_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_count_1_cry_1_c_LC_7_1_0 (
            .in0(_gnd_net_),
            .in1(N__903),
            .in2(N__802),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_1_0_),
            .carryout(un2_count_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_2_LC_7_1_1.C_ON=1'b1;
    defparam count_2_LC_7_1_1.SEQ_MODE=4'b1000;
    defparam count_2_LC_7_1_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_2_LC_7_1_1 (
            .in0(_gnd_net_),
            .in1(N__688),
            .in2(_gnd_net_),
            .in3(N__682),
            .lcout(countZ0Z_2),
            .ltout(),
            .carryin(un2_count_1_cry_1),
            .carryout(un2_count_1_cry_2),
            .clk(N__1154),
            .ce(),
            .sr(_gnd_net_));
    defparam count_3_LC_7_1_2.C_ON=1'b1;
    defparam count_3_LC_7_1_2.SEQ_MODE=4'b1000;
    defparam count_3_LC_7_1_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_3_LC_7_1_2 (
            .in0(_gnd_net_),
            .in1(N__679),
            .in2(_gnd_net_),
            .in3(N__673),
            .lcout(countZ0Z_3),
            .ltout(),
            .carryin(un2_count_1_cry_2),
            .carryout(un2_count_1_cry_3),
            .clk(N__1154),
            .ce(),
            .sr(_gnd_net_));
    defparam count_4_LC_7_1_3.C_ON=1'b1;
    defparam count_4_LC_7_1_3.SEQ_MODE=4'b1000;
    defparam count_4_LC_7_1_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_4_LC_7_1_3 (
            .in0(_gnd_net_),
            .in1(N__670),
            .in2(_gnd_net_),
            .in3(N__664),
            .lcout(countZ0Z_4),
            .ltout(),
            .carryin(un2_count_1_cry_3),
            .carryout(un2_count_1_cry_4),
            .clk(N__1154),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_5_LC_7_1_4.C_ON=1'b1;
    defparam count_RNO_0_5_LC_7_1_4.SEQ_MODE=4'b0000;
    defparam count_RNO_0_5_LC_7_1_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_5_LC_7_1_4 (
            .in0(_gnd_net_),
            .in1(N__819),
            .in2(_gnd_net_),
            .in3(N__736),
            .lcout(count_RNO_0Z0Z_5),
            .ltout(),
            .carryin(un2_count_1_cry_4),
            .carryout(un2_count_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_6_LC_7_1_5.C_ON=1'b1;
    defparam count_RNO_0_6_LC_7_1_5.SEQ_MODE=4'b0000;
    defparam count_RNO_0_6_LC_7_1_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 count_RNO_0_6_LC_7_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__778),
            .in3(N__733),
            .lcout(count_RNO_0Z0Z_6),
            .ltout(),
            .carryin(un2_count_1_cry_5),
            .carryout(un2_count_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_7_LC_7_1_6.C_ON=1'b1;
    defparam count_RNO_0_7_LC_7_1_6.SEQ_MODE=4'b0000;
    defparam count_RNO_0_7_LC_7_1_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_7_LC_7_1_6 (
            .in0(_gnd_net_),
            .in1(N__834),
            .in2(_gnd_net_),
            .in3(N__730),
            .lcout(count_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un2_count_1_cry_6),
            .carryout(un2_count_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_8_LC_7_1_7.C_ON=1'b1;
    defparam count_8_LC_7_1_7.SEQ_MODE=4'b1000;
    defparam count_8_LC_7_1_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_8_LC_7_1_7 (
            .in0(_gnd_net_),
            .in1(N__873),
            .in2(_gnd_net_),
            .in3(N__727),
            .lcout(countZ0Z_8),
            .ltout(),
            .carryin(un2_count_1_cry_7),
            .carryout(un2_count_1_cry_8),
            .clk(N__1154),
            .ce(),
            .sr(_gnd_net_));
    defparam count_9_LC_7_2_0.C_ON=1'b1;
    defparam count_9_LC_7_2_0.SEQ_MODE=4'b1000;
    defparam count_9_LC_7_2_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_9_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(N__885),
            .in2(_gnd_net_),
            .in3(N__724),
            .lcout(countZ0Z_9),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(un2_count_1_cry_9),
            .clk(N__1156),
            .ce(),
            .sr(_gnd_net_));
    defparam count_10_LC_7_2_1.C_ON=1'b1;
    defparam count_10_LC_7_2_1.SEQ_MODE=4'b1000;
    defparam count_10_LC_7_2_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_10_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(N__858),
            .in2(_gnd_net_),
            .in3(N__721),
            .lcout(countZ0Z_10),
            .ltout(),
            .carryin(un2_count_1_cry_9),
            .carryout(un2_count_1_cry_10),
            .clk(N__1156),
            .ce(),
            .sr(_gnd_net_));
    defparam count_11_LC_7_2_2.C_ON=1'b1;
    defparam count_11_LC_7_2_2.SEQ_MODE=4'b1000;
    defparam count_11_LC_7_2_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_11_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(N__847),
            .in2(_gnd_net_),
            .in3(N__718),
            .lcout(countZ0Z_11),
            .ltout(),
            .carryin(un2_count_1_cry_10),
            .carryout(un2_count_1_cry_11),
            .clk(N__1156),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_12_LC_7_2_3.C_ON=1'b1;
    defparam count_RNO_0_12_LC_7_2_3.SEQ_MODE=4'b0000;
    defparam count_RNO_0_12_LC_7_2_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_12_LC_7_2_3 (
            .in0(_gnd_net_),
            .in1(N__1045),
            .in2(_gnd_net_),
            .in3(N__715),
            .lcout(count_RNO_0Z0Z_12),
            .ltout(),
            .carryin(un2_count_1_cry_11),
            .carryout(un2_count_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_13_LC_7_2_4.C_ON=1'b1;
    defparam count_RNO_0_13_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam count_RNO_0_13_LC_7_2_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_13_LC_7_2_4 (
            .in0(_gnd_net_),
            .in1(N__1099),
            .in2(_gnd_net_),
            .in3(N__712),
            .lcout(count_RNO_0Z0Z_13),
            .ltout(),
            .carryin(un2_count_1_cry_12),
            .carryout(un2_count_1_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_14_LC_7_2_5.C_ON=1'b1;
    defparam count_RNO_0_14_LC_7_2_5.SEQ_MODE=4'b0000;
    defparam count_RNO_0_14_LC_7_2_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_14_LC_7_2_5 (
            .in0(_gnd_net_),
            .in1(N__1123),
            .in2(_gnd_net_),
            .in3(N__763),
            .lcout(count_RNO_0Z0Z_14),
            .ltout(),
            .carryin(un2_count_1_cry_13),
            .carryout(un2_count_1_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_15_LC_7_2_6.C_ON=1'b1;
    defparam count_15_LC_7_2_6.SEQ_MODE=4'b1000;
    defparam count_15_LC_7_2_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_15_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(N__940),
            .in2(_gnd_net_),
            .in3(N__760),
            .lcout(countZ0Z_15),
            .ltout(),
            .carryin(un2_count_1_cry_14),
            .carryout(un2_count_1_cry_15),
            .clk(N__1156),
            .ce(),
            .sr(_gnd_net_));
    defparam count_16_LC_7_2_7.C_ON=1'b1;
    defparam count_16_LC_7_2_7.SEQ_MODE=4'b1000;
    defparam count_16_LC_7_2_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_16_LC_7_2_7 (
            .in0(_gnd_net_),
            .in1(N__961),
            .in2(_gnd_net_),
            .in3(N__757),
            .lcout(countZ0Z_16),
            .ltout(),
            .carryin(un2_count_1_cry_15),
            .carryout(un2_count_1_cry_16),
            .clk(N__1156),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_17_LC_7_3_0.C_ON=1'b1;
    defparam count_RNO_0_17_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam count_RNO_0_17_LC_7_3_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_17_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__1066),
            .in2(_gnd_net_),
            .in3(N__754),
            .lcout(count_RNO_0Z0Z_17),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(un2_count_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_18_LC_7_3_1.C_ON=1'b1;
    defparam count_18_LC_7_3_1.SEQ_MODE=4'b1000;
    defparam count_18_LC_7_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_18_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__1441),
            .in2(_gnd_net_),
            .in3(N__751),
            .lcout(countZ0Z_18),
            .ltout(),
            .carryin(un2_count_1_cry_17),
            .carryout(un2_count_1_cry_18),
            .clk(N__1161),
            .ce(),
            .sr(_gnd_net_));
    defparam count_19_LC_7_3_2.C_ON=1'b1;
    defparam count_19_LC_7_3_2.SEQ_MODE=4'b1000;
    defparam count_19_LC_7_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_19_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(N__1418),
            .in2(_gnd_net_),
            .in3(N__748),
            .lcout(countZ0Z_19),
            .ltout(),
            .carryin(un2_count_1_cry_18),
            .carryout(un2_count_1_cry_19),
            .clk(N__1161),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_20_LC_7_3_3.C_ON=1'b1;
    defparam count_RNO_0_20_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam count_RNO_0_20_LC_7_3_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_20_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(N__1309),
            .in2(_gnd_net_),
            .in3(N__745),
            .lcout(count_RNO_0Z0Z_20),
            .ltout(),
            .carryin(un2_count_1_cry_19),
            .carryout(un2_count_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_21_LC_7_3_4.C_ON=1'b1;
    defparam count_RNO_0_21_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam count_RNO_0_21_LC_7_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 count_RNO_0_21_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__1321),
            .in2(_gnd_net_),
            .in3(N__742),
            .lcout(count_RNO_0Z0Z_21),
            .ltout(),
            .carryin(un2_count_1_cry_20),
            .carryout(un2_count_1_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_22_LC_7_3_5.C_ON=1'b0;
    defparam count_22_LC_7_3_5.SEQ_MODE=4'b1000;
    defparam count_22_LC_7_3_5.LUT_INIT=16'b0010001010001000;
    LogicCell40 count_22_LC_7_3_5 (
            .in0(N__1003),
            .in1(N__1333),
            .in2(_gnd_net_),
            .in3(N__739),
            .lcout(countZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1161),
            .ce(),
            .sr(_gnd_net_));
    defparam count_7_LC_8_1_0.C_ON=1'b0;
    defparam count_7_LC_8_1_0.SEQ_MODE=4'b1000;
    defparam count_7_LC_8_1_0.LUT_INIT=16'b1000000011001100;
    LogicCell40 count_7_LC_8_1_0 (
            .in0(N__1288),
            .in1(N__910),
            .in2(N__1216),
            .in3(N__1256),
            .lcout(countZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(_gnd_net_));
    defparam count_1_LC_8_1_1.C_ON=1'b0;
    defparam count_1_LC_8_1_1.SEQ_MODE=4'b1000;
    defparam count_1_LC_8_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 count_1_LC_8_1_1 (
            .in0(_gnd_net_),
            .in1(N__800),
            .in2(_gnd_net_),
            .in3(N__904),
            .lcout(countZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(_gnd_net_));
    defparam count_5_LC_8_1_2.C_ON=1'b0;
    defparam count_5_LC_8_1_2.SEQ_MODE=4'b1000;
    defparam count_5_LC_8_1_2.LUT_INIT=16'b1000000011001100;
    LogicCell40 count_5_LC_8_1_2 (
            .in0(N__1286),
            .in1(N__892),
            .in2(N__1215),
            .in3(N__1255),
            .lcout(countZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIOBUR_8_LC_8_1_3.C_ON=1'b0;
    defparam count_RNIOBUR_8_LC_8_1_3.SEQ_MODE=4'b0000;
    defparam count_RNIOBUR_8_LC_8_1_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 count_RNIOBUR_8_LC_8_1_3 (
            .in0(N__886),
            .in1(N__874),
            .in2(N__862),
            .in3(N__846),
            .lcout(),
            .ltout(op_lt_op_lt_count8lto11_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNITTD11_5_LC_8_1_4.C_ON=1'b0;
    defparam count_RNITTD11_5_LC_8_1_4.SEQ_MODE=4'b0000;
    defparam count_RNITTD11_5_LC_8_1_4.LUT_INIT=16'b0111000011110000;
    LogicCell40 count_RNITTD11_5_LC_8_1_4 (
            .in0(N__835),
            .in1(N__777),
            .in2(N__823),
            .in3(N__820),
            .lcout(op_lt_op_lt_count8lt14),
            .ltout(op_lt_op_lt_count8lt14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNICTR52_12_LC_8_1_5.C_ON=1'b0;
    defparam count_RNICTR52_12_LC_8_1_5.SEQ_MODE=4'b0000;
    defparam count_RNICTR52_12_LC_8_1_5.LUT_INIT=16'b1111011111111111;
    LogicCell40 count_RNICTR52_12_LC_8_1_5 (
            .in0(N__1129),
            .in1(N__1102),
            .in2(N__808),
            .in3(N__1048),
            .lcout(op_lt_op_lt_count8lto19_1_N_5),
            .ltout(op_lt_op_lt_count8lto19_1_N_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_0_LC_8_1_6.C_ON=1'b0;
    defparam count_0_LC_8_1_6.SEQ_MODE=4'b1000;
    defparam count_0_LC_8_1_6.LUT_INIT=16'b0101000100010001;
    LogicCell40 count_0_LC_8_1_6 (
            .in0(N__801),
            .in1(N__1254),
            .in2(N__805),
            .in3(N__1277),
            .lcout(countZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(_gnd_net_));
    defparam count_6_LC_8_1_7.C_ON=1'b0;
    defparam count_6_LC_8_1_7.SEQ_MODE=4'b1000;
    defparam count_6_LC_8_1_7.LUT_INIT=16'b1101010100000000;
    LogicCell40 count_6_LC_8_1_7 (
            .in0(N__1253),
            .in1(N__1287),
            .in2(N__1214),
            .in3(N__784),
            .lcout(countZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_1_22_LC_8_2_0.C_ON=1'b0;
    defparam count_RNO_1_22_LC_8_2_0.SEQ_MODE=4'b0000;
    defparam count_RNO_1_22_LC_8_2_0.LUT_INIT=16'b0001111100000000;
    LogicCell40 count_RNO_1_22_LC_8_2_0 (
            .in0(N__962),
            .in1(N__941),
            .in2(N__1076),
            .in3(N__1385),
            .lcout(),
            .ltout(op_lt_op_lt_count8lto22_2_0_tz_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_0_22_LC_8_2_1.C_ON=1'b0;
    defparam count_RNO_0_22_LC_8_2_1.SEQ_MODE=4'b0000;
    defparam count_RNO_0_22_LC_8_2_1.LUT_INIT=16'b1111010101110101;
    LogicCell40 count_RNO_0_22_LC_8_2_1 (
            .in0(N__1296),
            .in1(N__1024),
            .in2(N__1006),
            .in3(N__982),
            .lcout(count_RNO_0Z0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIAEV82_17_LC_8_2_2.C_ON=1'b0;
    defparam count_RNIAEV82_17_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam count_RNIAEV82_17_LC_8_2_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 count_RNIAEV82_17_LC_8_2_2 (
            .in0(N__1443),
            .in1(N__1297),
            .in2(N__1077),
            .in3(N__1419),
            .lcout(op_lt_op_lt_count8lto22),
            .ltout(op_lt_op_lt_count8lto22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_13_LC_8_2_3.C_ON=1'b0;
    defparam count_13_LC_8_2_3.SEQ_MODE=4'b1000;
    defparam count_13_LC_8_2_3.LUT_INIT=16'b1000110000001100;
    LogicCell40 count_13_LC_8_2_3 (
            .in0(N__1386),
            .in1(N__997),
            .in2(N__988),
            .in3(N__1364),
            .lcout(countZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1155),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIFVD41_12_LC_8_2_4.C_ON=1'b0;
    defparam count_RNIFVD41_12_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam count_RNIFVD41_12_LC_8_2_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 count_RNIFVD41_12_LC_8_2_4 (
            .in0(N__1047),
            .in1(N__1101),
            .in2(_gnd_net_),
            .in3(N__1125),
            .lcout(),
            .ltout(op_lt_op_lt_count8lto14_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNIRC5U2_15_LC_8_2_5.C_ON=1'b0;
    defparam count_RNIRC5U2_15_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam count_RNIRC5U2_15_LC_8_2_5.LUT_INIT=16'b0001000100000001;
    LogicCell40 count_RNIRC5U2_15_LC_8_2_5 (
            .in0(N__942),
            .in1(N__963),
            .in2(N__985),
            .in3(N__981),
            .lcout(op_lt_op_lt_count8lt17),
            .ltout(op_lt_op_lt_count8lt17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_12_LC_8_2_6.C_ON=1'b0;
    defparam count_12_LC_8_2_6.SEQ_MODE=4'b1000;
    defparam count_12_LC_8_2_6.LUT_INIT=16'b1100010001000100;
    LogicCell40 count_12_LC_8_2_6 (
            .in0(N__1252),
            .in1(N__973),
            .in2(N__967),
            .in3(N__1387),
            .lcout(countZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1155),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNI45JG1_15_LC_8_2_7.C_ON=1'b0;
    defparam count_RNI45JG1_15_LC_8_2_7.SEQ_MODE=4'b0000;
    defparam count_RNI45JG1_15_LC_8_2_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 count_RNI45JG1_15_LC_8_2_7 (
            .in0(N__1420),
            .in1(N__964),
            .in2(N__946),
            .in3(N__1442),
            .lcout(op_lt_op_lt_count8lto19_1_m4_i_a3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_21_LC_8_3_0.C_ON=1'b0;
    defparam count_21_LC_8_3_0.SEQ_MODE=4'b1000;
    defparam count_21_LC_8_3_0.LUT_INIT=16'b1011001100000000;
    LogicCell40 count_21_LC_8_3_0 (
            .in0(N__1389),
            .in1(N__1261),
            .in2(N__1366),
            .in3(N__925),
            .lcout(countZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1157),
            .ce(),
            .sr(_gnd_net_));
    defparam count_17_LC_8_3_3.C_ON=1'b0;
    defparam count_17_LC_8_3_3.SEQ_MODE=4'b1000;
    defparam count_17_LC_8_3_3.LUT_INIT=16'b1101000001010000;
    LogicCell40 count_17_LC_8_3_3 (
            .in0(N__1259),
            .in1(N__1363),
            .in2(N__919),
            .in3(N__1390),
            .lcout(countZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1157),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNILL9O_18_LC_8_3_4.C_ON=1'b0;
    defparam count_RNILL9O_18_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam count_RNILL9O_18_LC_8_3_4.LUT_INIT=16'b0000000000001111;
    LogicCell40 count_RNILL9O_18_LC_8_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1444),
            .in3(N__1417),
            .lcout(op_lt_op_lt_count8lto19_0),
            .ltout(op_lt_op_lt_count8lto19_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam count_14_LC_8_3_5.C_ON=1'b0;
    defparam count_14_LC_8_3_5.SEQ_MODE=4'b1000;
    defparam count_14_LC_8_3_5.LUT_INIT=16'b1100010001000100;
    LogicCell40 count_14_LC_8_3_5 (
            .in0(N__1258),
            .in1(N__1399),
            .in2(N__1393),
            .in3(N__1362),
            .lcout(countZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1157),
            .ce(),
            .sr(_gnd_net_));
    defparam count_20_LC_8_3_6.C_ON=1'b0;
    defparam count_20_LC_8_3_6.SEQ_MODE=4'b1000;
    defparam count_20_LC_8_3_6.LUT_INIT=16'b1011001100000000;
    LogicCell40 count_20_LC_8_3_6 (
            .in0(N__1388),
            .in1(N__1260),
            .in2(N__1365),
            .in3(N__1339),
            .lcout(countZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1157),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNICVG41_22_LC_8_3_7.C_ON=1'b0;
    defparam count_RNICVG41_22_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam count_RNICVG41_22_LC_8_3_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 count_RNICVG41_22_LC_8_3_7 (
            .in0(N__1332),
            .in1(N__1320),
            .in2(_gnd_net_),
            .in3(N__1308),
            .lcout(op_lt_op_lt_count8lto22_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ledZ0_LC_9_1_1.C_ON=1'b0;
    defparam ledZ0_LC_9_1_1.SEQ_MODE=4'b1000;
    defparam ledZ0_LC_9_1_1.LUT_INIT=16'b1011010000111100;
    LogicCell40 ledZ0_LC_9_1_1 (
            .in0(N__1285),
            .in1(N__1257),
            .in2(N__1182),
            .in3(N__1213),
            .lcout(led_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1152),
            .ce(),
            .sr(_gnd_net_));
    defparam count_RNO_2_22_LC_9_2_0.C_ON=1'b0;
    defparam count_RNO_2_22_LC_9_2_0.SEQ_MODE=4'b0000;
    defparam count_RNO_2_22_LC_9_2_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 count_RNO_2_22_LC_9_2_0 (
            .in0(N__1124),
            .in1(N__1100),
            .in2(N__1078),
            .in3(N__1046),
            .lcout(op_lt_op_lt_count8lto22_d_a0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_30_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_30_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // Blink
