Blinky_pll_inst: Blinky_pll
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
