Blinky_pll_inst: Blinky_pll
port map(
          REFERENCECLK => REFERENCECLK ,
          PLLOUTCORE =>PLLOUTCORE ,
          PLLOUTGLOBAL =>PLLOUTGLOBAL ,
          RESET =>RESET 
        );
